module ksa(cy,s,a,b,cin);
input [7:0]a,b;
input cin;
output [7:0]s;
output cy;
wire [7:0]p,g;
wire [7:0]c,g1,g2,g3;
assign p[0]=a[0]^b[0];
assign p[1]=a[1]^b[1];
assign p[2]=a[2]^b[2];
assign p[3]=a[3]^b[3];
assign p[4]=a[4]^b[4];
assign p[5]=a[5]^b[5];
assign p[6]=a[6]^b[6];
assign p[7]=a[7]^b[7];
assign g[0]=a[0]&b[0];
assign g[1]=a[1]&b[1];
assign g[2]=a[2]&b[2];
assign g[3]=a[3]&b[3];
assign g[4]=a[4]&b[4];
assign g[5]=a[5]&b[5];
assign g[6]=a[6]&b[6];
assign g[7]=a[7]&b[7];
assign g1[0]=g[0];
assign g1[1]=g[1]|(p[0]&g[0]);
assign g1[2]=g[2]|(p[1]&g[1]);
assign g1[3]=g[3]|(p[2]&g[2]);
assign g1[4]=g[4]|(p[3]&g[3]);
assign g1[5]=g[5]|(p[4]&g[4]);
assign g1[6]=g[6]|(p[5]&g[5]);
assign g1[7]=g[7]|(p[6]&g[6]);
assign g2[0]=g1[0];
assign g2[1]=g1[1];
assign g2[2]=g1[2]|(p[0]&g1[0]);
assign g2[3]=g1[3]|(p[1]&g2[1]);
assign g2[4]=g2[4] |(p[2]&g2[2]);
assign g2[5]=g2[5] |(p[3]&g2[3]);
assign g2[6]=g2[6] |(p[4]&g2[4]);
assign g2[7]=g2[7] |(p[5]&g2[5]);
assign g3[0]=g1[0];
assign g3[1]=g1[1];
assign g3[2]=g1[2];
assign g3[3]=g1[3];
assign g3[4]=g2[4] |(p[0]&g2[2]);
assign g3[5]=g2[5] |(p[1]&g2[3]);
assign g3[6]=g2[6] |(p[2]&g2[4]);
assign g3[7]=g2[7] |(p[3]&g2[3]);
assign c[0]=cin;
assign c[1]=g[0]|(p[0]&cin);
assign c[2]=g[1]|(p[1]&c[1]);
assign c[3]=g[2]|(p[2]&c[2]);
assign c[4]=g[3]|(p[3]&c[3]);
assign c[5]=g[4]|(p[4]&c[4]);
assign c[6]=g[5]|(p[5]&c[5]);
assign c[7]=g[6]|(p[6]&c[6]);
assign cy=g[7]|(p[7]&c[7]);
assign s[0]=p[0]^cin;
assign s[1]=p[1]^c[1];
assign s[2]=p[2]^c[2];
assign s[3]=p[3]^c[3];
assign s[4]=p[4]^c[4];
assign s[5]=p[5]^c[5];
assign s[6]=p[6]^c[6];
assign s[7]=p[7]^c[7];
endmodule
