module testbench;

reg [3:0]I;
wire [1:0]O;
priority_encoder uut(.I(I),.O(O));
initial begin
    I = 4'b0000; #10;
    I = 4'b0001; #10;
    I = 4'b0010; #10;
    I = 4'b0011; #10;
    I = 4'b0100; #10;
    I = 4'b0101; #10;
    I = 4'b0110; #10;
    I = 4'b0111; #10;
    I = 4'b1110; #10;
    I = 4'b1111; #10;
    
       
$finish;
end
endmodule
